*rc circuit with ac analysis
vcc in 0 AC 1
r1 in out 1k
c1 out 0 1u
.ac dec 100 1 100k
.end
