*voltage+current+resistor
v1 1 0 1
r1 1 2 1k
r2 2 0 2k
r3 2 3 3k
i1 0 3 1m
.op
.end
