*lcr circuit
vcc 1 0 ac 1
r1  1 2 6
l1  2 3 .0015923
c1  3 0 .000796178344
.ac dec 10 1 20k
.end
