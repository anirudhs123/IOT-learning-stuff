*voltage divider
V1 1 0 12
R1 1 2 2500
c1 2 0 1

.op
.end
