* forward bias led
V1 1 0 sin(0 1 1k)
R1 1 2 1k
*D1 2 0 LED2
*d2 2 0 led1
d3 2 0 led3
*Typ RED GaAs LED:  Vf=1.7V Vr If=40mA trr=3uS
*.MODEL LED1 D (IS=93.2P RS=42M N=3.73 BV=4 IBV=10U
*+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)
*Typ RED,GREEN,YELLOW,AMBER GaAs LED: Vf=2.1V Vr=4V If=40mA trr=3uS
*.MODEL LED2 D (IS=93.1P RS=42M N=4.61 BV=4 IBV=10U
*+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)

*Typ BLUE SiC LED: Vf=3.4V Vr=5V If=40mA trr=3uS
.MODEL LED3 D (IS=93.1P RS=42M N=7.47 BV=5 IBV=30U
+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)

*.lib C:\Users\dell\Documents\LTspiceXVII\lib\cmp\standard.dio
.tran 5m

.end
