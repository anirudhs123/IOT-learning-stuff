*rc circuit with unit step voltage source
vcc in 0 pwl(0 0  0.0001m 5 1m 5)
r1 in out 1k
c1 out 0 1u
.tran 10m
.end
