*lcr circuit
vcc 1 0 sin(0 10 1k)
r1  1 2 6
l1  2 3 .0015923
c1  3 0 .000796178344
.tran 10m
.end
