*full wave rectifier
vs in  0 0
r1 out 0 5k
d1 in out dmod
d2 out in dmod
.model dmod D(Is=153.4e-12 N=1.487 Rs=.6329 Ikf=3.53m Xti=3 Eg=1.11 cjo=2.51p
+           M=.1575 Vj=.5 Fc=.5 Isr=4.763n Nr=2 Bv=35 Ibv=5u Tt=5.771n)
.dc vs -2 2 1m
.end
